Series combination of two transistors
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.18u
.param width_P=20*LAMBDA
.param width_N=10*LAMBDA
.global gnd vdd

VDS D gnd 0
VGS G gnd 1.8V

M1 D G gnd gnd CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA}


.dc VDS 0 10 0.1


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
let x = (-VDS#branch)
set curplottitle="Id vs Vds Characteristics"
plot x 

hardcopy fig_Q4a.eps (-VDS#branch)
.endc