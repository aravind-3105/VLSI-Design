VLSI Assignment Question 6bii
* Answers to question 6b (ii)
.include TSMC_180nm.txt
.param SUPPLY=-1V
.param LAMBDA=0.09u
.param width_P=20*LAMBDA
.global gnd vdd

Vdd	 y gnd 0V
vin x gnd 0V

M1 x y z supply CMOSP W={width_P} L={2*LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

Cout z gnd 100f

.tran 0.001n 100n
.ic v(z)= 1.8
.ic v(y) = 1.8

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
*plot v(a)
*plot v(b)
plot  v(z)

hardcopy fig_Q6b_ii.eps v(z)
.endc




