magic
tech scmos
timestamp 1613681421
<< nwell >>
rect 0 0 24 37
<< ntransistor >>
rect 11 -18 13 -8
<< ptransistor >>
rect 11 6 13 31
<< ndiffusion >>
rect 10 -18 11 -8
rect 13 -18 14 -8
<< pdiffusion >>
rect 10 6 11 31
rect 13 6 14 31
<< ndcontact >>
rect 6 -18 10 -8
rect 14 -18 18 -8
<< pdcontact >>
rect 6 6 10 31
rect 14 6 18 31
<< polysilicon >>
rect 11 31 13 34
rect 11 -8 13 6
rect 11 -28 13 -18
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 0 35 24 39
rect 6 31 10 35
rect 14 -1 18 6
rect 0 -5 7 -1
rect 14 -5 24 -1
rect 14 -8 18 -5
rect 6 -29 10 -18
rect 0 -33 24 -29
<< end >>
