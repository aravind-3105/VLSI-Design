.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
vin_x x 0 pulse 0 1.8 0ns 100ps 100ps 4.9ns 10ns

.subckt inv yi xi vdd gnd
M1      yi       xi       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      yi       xi       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

.subckt MUX2_1 x x_bar y vdd gnd 
    M1      vdd       x       y     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    M2      y         x_bar   gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}     
.ends MUX2_1


x0 x_bar x vdd gnd inv
x1 x x_bar y vdd gnd MUX2_1


.tran 0.1n 100n

.control
* set hcopypscolor = 1
* set color0=white
* set color1=black

run
plot v(x) v(x_bar) v(y) 
plot v(x_bar) 
plot v(y) 
set curplottitle= "Aravind Narayanan-2019102014"
.endc
