magic
tech scmos
timestamp 1613808346
<< metal1 >>
rect -27 68 360 73
rect -27 -68 -20 68
rect -16 28 4 32
rect 14 28 31 32
rect 38 28 55 32
rect 62 28 79 32
rect 86 28 103 32
rect 110 28 127 32
rect 134 28 151 32
rect 158 28 175 32
rect 182 28 199 32
rect 206 28 223 32
rect 230 28 247 32
rect 254 28 271 32
rect 278 28 295 32
rect 302 28 319 32
rect 326 28 343 32
rect 350 28 394 32
rect -16 -40 -9 28
rect -1 -4 384 4
rect 389 -40 394 28
rect -16 -44 10 -40
rect 17 -44 34 -40
rect 41 -44 58 -40
rect 65 -44 82 -40
rect 89 -44 106 -40
rect 113 -44 130 -40
rect 137 -44 154 -40
rect 161 -44 178 -40
rect 185 -44 202 -40
rect 209 -44 226 -40
rect 233 -44 250 -40
rect 257 -44 274 -40
rect 281 -44 298 -40
rect 305 -44 322 -40
rect 329 -44 346 -40
rect 353 -44 370 -40
rect 384 -44 394 -40
rect -27 -72 2 -68
use inverter_wo_label_Q5  inverter_wo_label_Q5_0
array 0 14 24 0 0 72
timestamp 1613681421
transform 1 0 0 0 1 33
box 0 -33 24 39
use inverter_wo_label_Q5  inverter_wo_label_Q5_1
array 0 15 -24 0 0 72
timestamp 1613681421
transform -1 0 24 0 1 -39
box 0 -33 24 39
<< labels >>
rlabel metal1 0 68 360 73 5 vdd
rlabel metal1 -1 -4 384 4 1 gnd
rlabel metal1 -16 28 4 32 1 M1
rlabel metal1 14 28 31 32 1 M2
rlabel metal1 38 28 55 32 1 M3
rlabel metal1 62 28 79 32 1 M4
rlabel metal1 86 28 103 32 1 M5
rlabel metal1 110 28 127 32 1 M6
rlabel metal1 134 28 151 32 1 M7
rlabel metal1 158 28 175 32 1 M8
rlabel metal1 182 28 199 32 1 M9
rlabel metal1 206 28 223 32 1 M10
rlabel metal1 230 28 247 32 1 M11
rlabel metal1 254 28 271 32 1 M12
rlabel metal1 278 28 295 32 1 M13
rlabel metal1 302 28 319 32 1 M14
rlabel metal1 326 28 343 32 1 M15
rlabel metal1 350 28 393 32 1 M16
rlabel metal1 353 -44 370 -40 1 M17
rlabel metal1 329 -44 346 -40 1 M18
rlabel metal1 305 -44 322 -40 1 M19
rlabel metal1 281 -44 298 -40 1 M20
rlabel metal1 257 -44 274 -40 1 M21
rlabel metal1 233 -44 250 -40 1 M22
rlabel metal1 209 -44 226 -40 1 M23
rlabel metal1 185 -44 202 -40 1 M24
rlabel metal1 161 -44 178 -40 1 M25
rlabel metal1 137 -44 154 -40 1 M26
rlabel metal1 113 -44 130 -40 1 M27
rlabel metal1 89 -44 106 -40 1 M28
rlabel metal1 65 -44 82 -40 1 M29
rlabel metal1 41 -44 58 -40 1 M30
rlabel metal1 17 -44 34 -40 1 M31
<< end >>
