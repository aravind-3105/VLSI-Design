.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={2.5*width_N}
.global gnd vdd

.subckt inv y x vdd gnd
M1      y       x       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      y       x       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

x1 1 in vdd gnd inv
x2 2 1 vdd gnd inv
x3 3 2 vdd gnd inv
x4 4 3 vdd gnd inv
x5 5 4 vdd gnd inv
x6 6 5 vdd gnd inv
x7 7 6 vdd gnd inv
x8 8 7 vdd gnd inv
x9 9 8 vdd gnd inv
x10 10 9 vdd gnd inv
x11 11 10 vdd gnd inv
x12 12 11 vdd gnd inv
x13 13 12 vdd gnd inv
x14 14 13 vdd gnd inv
x15 15 14 vdd gnd inv
x16 16 15 vdd gnd inv
x17 17 16 vdd gnd inv
x18 18 17 vdd gnd inv
x19 19 18 vdd gnd inv
x20 20 19 vdd gnd inv
x21 21 20 vdd gnd inv
x22 22 21 vdd gnd inv
x23 23 22 vdd gnd inv
x24 24 23 vdd gnd inv
x25 25 24 vdd gnd inv
x26 26 25 vdd gnd inv
x27 27 26 vdd gnd inv
x28 28 27 vdd gnd inv
x29 29 28 vdd gnd inv
x30 30 29 vdd gnd inv
x31 in 30 vdd gnd inv

Vdd	vdd	gnd	'SUPPLY'

.ic v(in) = 'SUPPLY'
.tran 10n 20n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
set curplottitle="v(out)"
plot v(in)

.endc