* SPICE3 file created from new1_optimized_ring_oscillator.ext - technology: scmos

.option scale=0.09u

M1000 M1 M31 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=3875 ps=1860
M1001 M1 M31 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=1550 ps=930
M1002 M31 M30 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1003 M31 M30 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 M30 M29 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1005 M30 M29 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1006 M29 M28 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1007 M29 M28 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1008 M28 M27 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1009 M28 M27 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1010 M27 M26 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1011 M27 M26 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1012 M26 M25 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1013 M26 M25 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 M25 M24 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1015 M25 M24 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 M24 M23 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1017 M24 M23 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1018 M23 M22 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1019 M23 M22 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1020 M22 M21 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1021 M22 M21 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1022 M21 M20 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1023 M21 M20 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1024 M20 M19 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1025 M20 M19 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 M19 M18 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1027 M19 M18 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1028 M18 M17 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1029 M18 M17 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1030 M17 M16 vdd inverter_wo_label_Q5_1[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1031 M17 M16 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1032 M2 M1 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1033 M2 M1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1034 M3 M2 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1035 M3 M2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1036 M4 M3 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1037 M4 M3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 M5 M4 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1039 M5 M4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 M6 M5 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1041 M6 M5 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1042 M7 M6 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1043 M7 M6 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1044 M8 M7 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1045 M8 M7 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1046 M9 M8 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1047 M9 M8 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1048 M10 M9 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1049 M10 M9 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 M11 M10 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1051 M11 M10 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1052 M12 M11 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1053 M12 M11 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1054 M13 M12 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1055 M13 M12 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1056 M14 M13 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1057 M14 M13 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1058 M15 M14 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1059 M15 M14 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 M16 M15 vdd inverter_wo_label_Q5_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1061 M16 M15 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 inverter_wo_label_Q5_1[0]/w_0_0# vdd 1.2fF
C1 vdd M1 1.2fF
C2 inverter_wo_label_Q5_0[0]/w_0_0# vdd 1.2fF
C3 vdd gnd! 1.9fF
C4 inverter_wo_label_Q5_0[0]/w_0_0# gnd! 13.4fF
C5 gnd gnd! 3.2fF
C6 M16 gnd! 1.3fF
C7 inverter_wo_label_Q5_1[0]/w_0_0# gnd! 14.3fF
C8 M30 gnd! 1.1fF
C9 M31 gnd! 1.2fF
C10 M1 gnd! 2.3fF
