magic
tech scmos
timestamp 1613672100
<< metal1 >>
rect 0 99 75 102
rect -9 33 2 37
rect 14 33 30 37
rect 39 33 55 37
rect 75 33 85 37
rect -9 -5 -4 33
rect 0 0 75 3
rect 80 -5 85 33
rect -9 -8 85 -5
use inverter  inverter_0
array 0 2 25 0 0 101
timestamp 1613670903
transform 1 0 9 0 1 38
box -9 -38 16 64
<< labels >>
rlabel metal1 0 0 75 0 1 gnd
rlabel metal1 0 102 75 102 5 vdd
rlabel metal1 -9 -8 85 -5 1 m1
rlabel metal1 14 33 30 37 1 m2
rlabel metal1 39 33 55 37 1 m3
<< end >>
