* SPICE3 file created from ro2.ext - technology: scmos

.option scale=0.09u

M1000 basicinv_0[1]/a_7_n5# 16 vdd basicinv_0[0]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=3875 ps=1860
M1001 basicinv_0[1]/a_7_n5# 16 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=1550 ps=930
M1002 basicinv_0[2]/a_7_n5# basicinv_0[1]/a_7_n5# vdd basicinv_0[1]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1003 basicinv_0[2]/a_7_n5# basicinv_0[1]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 basicinv_0[3]/a_7_n5# basicinv_0[2]/a_7_n5# vdd basicinv_0[2]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1005 basicinv_0[3]/a_7_n5# basicinv_0[2]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1006 basicinv_0[4]/a_7_n5# basicinv_0[3]/a_7_n5# vdd basicinv_0[3]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1007 basicinv_0[4]/a_7_n5# basicinv_0[3]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1008 basicinv_0[5]/a_7_n5# basicinv_0[4]/a_7_n5# vdd basicinv_0[4]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1009 basicinv_0[5]/a_7_n5# basicinv_0[4]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1010 basicinv_0[6]/a_7_n5# basicinv_0[5]/a_7_n5# vdd basicinv_0[5]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1011 basicinv_0[6]/a_7_n5# basicinv_0[5]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1012 basicinv_0[7]/a_7_n5# basicinv_0[6]/a_7_n5# vdd basicinv_0[6]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1013 basicinv_0[7]/a_7_n5# basicinv_0[6]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 basicinv_0[8]/a_7_n5# basicinv_0[7]/a_7_n5# vdd basicinv_0[7]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1015 basicinv_0[8]/a_7_n5# basicinv_0[7]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 basicinv_0[9]/a_7_n5# basicinv_0[8]/a_7_n5# vdd basicinv_0[8]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1017 basicinv_0[9]/a_7_n5# basicinv_0[8]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1018 basicinv_0[10]/a_7_n5# basicinv_0[9]/a_7_n5# vdd basicinv_0[9]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1019 basicinv_0[10]/a_7_n5# basicinv_0[9]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1020 basicinv_0[11]/a_7_n5# basicinv_0[10]/a_7_n5# vdd basicinv_0[10]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1021 basicinv_0[11]/a_7_n5# basicinv_0[10]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1022 basicinv_0[12]/a_7_n5# basicinv_0[11]/a_7_n5# vdd basicinv_0[11]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1023 basicinv_0[12]/a_7_n5# basicinv_0[11]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1024 basicinv_0[13]/a_7_n5# basicinv_0[12]/a_7_n5# vdd basicinv_0[12]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1025 basicinv_0[13]/a_7_n5# basicinv_0[12]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 basicinv_0[14]/a_7_n5# basicinv_0[13]/a_7_n5# vdd basicinv_0[13]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1027 basicinv_0[14]/a_7_n5# basicinv_0[13]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1028 in basicinv_0[14]/a_7_n5# vdd basicinv_0[14]/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1029 in basicinv_0[14]/a_7_n5# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1030 16 15 vdd basicinv_1/w_0_0# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1031 16 15 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1032 15 14 vdd w_2_423# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1033 15 14 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1034 14 13 vdd w_2_393# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1035 14 13 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1036 13 12 vdd w_2_363# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1037 13 12 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 12 11 vdd w_2_333# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1039 12 11 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 11 10 vdd w_2_303# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1041 11 10 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1042 10 9 vdd w_2_273# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1043 10 9 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1044 9 8 vdd w_2_243# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1045 9 8 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1046 8 7 vdd w_2_213# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1047 8 7 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1048 7 6 vdd w_2_183# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1049 7 6 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 6 5 vdd w_2_153# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1051 6 5 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1052 5 4 vdd w_2_123# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1053 5 4 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1054 4 3 vdd w_2_93# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1055 4 3 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1056 3 2 vdd w_2_63# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1057 3 2 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1058 2 1 vdd w_2_33# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1059 2 1 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 1 in vdd w_2_3# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1061 1 in gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 w_2_33# gnd! 1.0fF
C1 w_2_63# gnd! 1.0fF
C2 w_2_93# gnd! 1.0fF
C3 w_2_123# gnd! 1.0fF
C4 w_2_153# gnd! 1.0fF
C5 w_2_183# gnd! 1.0fF
C6 w_2_213# gnd! 1.0fF
C7 w_2_243# gnd! 1.0fF
C8 w_2_273# gnd! 1.0fF
C9 w_2_303# gnd! 1.0fF
C10 w_2_333# gnd! 1.0fF
C11 w_2_363# gnd! 1.0fF
C12 w_2_393# gnd! 1.0fF
C13 w_2_423# gnd! 1.0fF
C14 gnd gnd! 6.4fF
C15 basicinv_1/w_0_0# gnd! 1.0fF
C16 vdd gnd! 8.4fF