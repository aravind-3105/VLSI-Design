* SPICE3 file created from inverter.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
vin inp gnd pulse 0 1.8 0ns 1ns 1ns 10ns 20ns

.option scale=0.09u

M1000 x inp vdd w_n9_0# CMOSP w=50 l=2
+  ad=250 pd=110 as=500 ps=220

M1001 out x vdd w_n9_0# CMOSP w=50 l=2
+  ad=250 pd=110 as=0 ps=0

M1002 x inp gnd gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100

M1003 out x gnd gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0

C0 w_n9_0# gnd 2.8fF
*Cout out gnd 100f
.tran 0.01n 80n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))
run 
plot v(out) v(inp)
set hcopypscolor = 1
hardcopy Inverter_post.eps v(inp) v(out)
.endc
.end