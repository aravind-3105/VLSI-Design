* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.09u

M1000 output input vdd w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=250 ps=110
M1001 output input gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
C0 w_n9_0# gnd! 1.6fF
