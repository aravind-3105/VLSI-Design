* SPICE3 file created from double.ext - technology: scmos

.option scale=0.09u

M1000 mid in vdd w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=80 ps=52
M1001 out mid vdd w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1002 mid in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1003 out mid gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 w_0_0# gnd! 1.1fF
