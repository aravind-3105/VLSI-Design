VLSI Assignment Question 6aii
* Answers to question 6a (ii)
.include TSMC_180nm.txt
.param SUPPLY=-2.8V
.param LAMBDA=0.09u
.param width_P=20*LAMBDA
.global gnd vdd

Vdd	 vdd gnd 'SUPPLY'
vin x gnd 0V

M1 z vdd x x CMOSP W={width_P} L={2*LAMBDA} +
AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

Cout z gnd 100f

.ic v(z)= 1.8
.tran 0.001n 5n



.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
*plot v(a)
*plot v(b)
plot  v(z)

hardcopy fig_Q6b_ii.eps v(z)
.endc




