magic
tech scmos
timestamp 1613690691
<< metal1 >>
rect -24 68 360 74
rect -23 -68 -16 68
rect -8 28 3 32
rect 14 28 31 32
rect 38 28 55 32
rect 62 28 79 32
rect 86 28 103 32
rect 110 28 127 32
rect 134 28 151 32
rect 158 28 175 32
rect 182 28 199 32
rect 206 28 223 32
rect 230 28 247 32
rect 254 28 271 32
rect 278 28 295 32
rect 302 28 319 32
rect 326 28 343 32
rect 360 28 393 32
rect -8 -28 -4 28
rect 0 -4 384 4
rect 387 -28 393 28
rect -8 -32 7 -28
rect 14 -32 31 -28
rect 38 -32 55 -28
rect 62 -32 79 -28
rect 86 -32 103 -28
rect 110 -32 127 -28
rect 134 -32 151 -28
rect 158 -32 175 -28
rect 182 -32 199 -28
rect 206 -32 223 -28
rect 230 -32 247 -28
rect 254 -32 271 -28
rect 278 -32 295 -28
rect 302 -32 319 -28
rect 326 -32 343 -28
rect 350 -32 367 -28
rect 374 -32 393 -28
rect -23 -73 384 -68
use inverter_wo_label_Q5  inverter_wo_label_Q5_0
array 0 14 24 0 0 72
timestamp 1613681421
transform 1 0 0 0 1 33
box 0 -33 24 39
use inverter_wo_label_Q5  inverter_wo_label_Q5_1
array 0 15 24 0 0 -72
timestamp 1613681421
transform 1 0 0 0 -1 -33
box 0 -33 24 39
<< labels >>
rlabel metal1 -24 68 360 74 5 vdd
rlabel metal1 0 -4 384 4 1 gnd
rlabel metal1 14 28 31 32 1 M2
rlabel metal1 38 28 55 32 1 M3
rlabel metal1 62 28 79 32 1 M4
rlabel metal1 86 28 103 32 1 M5
rlabel metal1 110 28 127 32 1 M6
rlabel metal1 134 28 151 32 1 M7
rlabel metal1 158 28 175 32 1 M8
rlabel metal1 182 28 199 32 1 M9
rlabel metal1 206 28 223 32 1 M10
rlabel metal1 230 28 247 32 1 M11
rlabel metal1 254 28 271 32 1 M12
rlabel metal1 278 28 295 32 1 M13
rlabel metal1 302 28 319 32 1 M14
rlabel metal1 326 28 343 32 1 M15
rlabel metal1 326 -32 343 -28 1 M18
rlabel metal1 302 -32 319 -28 1 M19
rlabel metal1 158 -32 175 -28 1 M25
rlabel metal1 134 -32 151 -28 1 M26
rlabel metal1 110 -32 127 -28 1 M27
rlabel metal1 86 -32 103 -28 1 M28
rlabel metal1 62 -32 79 -28 1 M29
rlabel metal1 38 -32 55 -28 1 M30
rlabel metal1 14 -32 31 -28 1 M31
rlabel metal1 350 -32 367 -28 1 M17
rlabel metal1 278 -32 295 -28 1 M20
rlabel metal1 254 -32 271 -28 1 M21
rlabel metal1 230 -32 247 -28 1 M22
rlabel metal1 206 -32 223 -28 1 M23
rlabel metal1 182 -32 199 -28 1 M24
rlabel metal1 -8 28 3 32 1 M1
rlabel space 350 28 393 32 1 M16
<< end >>
