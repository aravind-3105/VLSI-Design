magic
tech scmos
timestamp 1613683967
<< metal1 >>
rect 0 68 744 73
rect -16 28 1 32
rect 14 28 31 32
rect 38 28 55 32
rect 62 28 79 32
rect 86 28 103 32
rect 110 28 127 32
rect 134 28 151 32
rect 158 28 175 32
rect 182 28 199 32
rect 206 28 223 32
rect 230 28 247 32
rect 254 28 271 32
rect 278 28 295 32
rect 302 28 319 32
rect 326 28 343 32
rect 350 28 367 32
rect 374 28 391 32
rect 398 28 415 32
rect 422 28 439 32
rect 446 28 463 32
rect 470 28 487 32
rect 494 28 511 32
rect 518 28 535 32
rect 566 28 583 32
rect 590 28 607 32
rect 614 28 631 32
rect 638 28 655 32
rect 662 28 679 32
rect 686 28 703 32
rect 710 28 727 32
rect 734 28 757 32
rect -16 -3 -8 28
rect 0 0 744 4
rect 751 -3 757 28
rect -16 -9 757 -3
use inverter_wo_label_Q5  inverter_wo_label_Q5_0
array 0 30 24 0 0 72
timestamp 1613681421
transform 1 0 0 0 1 33
box 0 -33 24 39
<< labels >>
rlabel metal1 0 0 744 4 1 gnd
rlabel metal1 0 68 744 73 5 vdd
rlabel metal1 14 28 31 32 1 M2
rlabel metal1 38 28 55 32 1 M3
rlabel metal1 62 28 79 32 1 M4
rlabel metal1 86 28 103 32 1 M5
rlabel metal1 110 28 127 32 1 M6
rlabel metal1 134 28 151 32 1 M7
rlabel metal1 158 28 175 32 1 M8
rlabel metal1 182 28 199 32 1 M9
rlabel metal1 206 28 223 32 1 M10
rlabel metal1 230 28 247 32 1 M11
rlabel metal1 254 28 271 32 1 M12
rlabel metal1 278 28 295 32 1 M13
rlabel metal1 302 28 319 32 1 M14
rlabel metal1 326 28 343 32 1 M15
rlabel metal1 350 28 367 32 1 M16
rlabel metal1 374 28 391 32 1 M17
rlabel metal1 398 28 415 32 1 M18
rlabel metal1 422 28 439 32 1 M19
rlabel metal1 446 28 463 32 1 M20
rlabel metal1 470 28 487 32 1 M21
rlabel metal1 494 28 511 32 1 M22
rlabel metal1 518 28 535 32 1 M23
rlabel space 542 28 559 32 1 M24
rlabel metal1 566 28 583 32 1 M25
rlabel metal1 590 28 607 32 1 M26
rlabel metal1 614 28 631 32 1 M27
rlabel metal1 638 28 655 32 1 M28
rlabel metal1 662 28 679 32 1 M29
rlabel metal1 686 28 703 32 1 M30
rlabel metal1 710 28 727 32 1 M31
rlabel metal1 734 28 757 32 1 M1
<< end >>
