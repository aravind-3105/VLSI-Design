.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={2.5*width_N}
.global gnd vdd

.option scale=0.09u

M1000 x in vdd w_n6_n6# CMOSP w=50 l=2
+  ad=250 pd=110 as=500 ps=220
M1001 out x vdd w_25_n6# CMOSP w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1002 x in gnd gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1003 out x gnd gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0

C0 w_25_n6# gnd 1.5fF
C1 w_n6_n6# gnd 1.5fF

Vdd	vdd	gnd	'SUPPLY'
vin in gnd 0

.dc vin 0 'SUPPLY' 0.01


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
set curplottitle="Vb vs Va"
plot v(x)

set curplottitle="d(Vb)/d(Va) vs Va"
plot deriv(v(x))/deriv(v(in))

.endc