magic
tech scmos
timestamp 1613668076
<< nwell >>
rect -9 0 16 63
<< ntransistor >>
rect 2 -30 4 -10
<< ptransistor >>
rect 2 6 4 56
<< ndiffusion >>
rect 1 -30 2 -10
rect 4 -30 5 -10
<< pdiffusion >>
rect 1 6 2 56
rect 4 6 5 56
<< ndcontact >>
rect -3 -30 1 -10
rect 5 -30 9 -10
<< pdcontact >>
rect -3 6 1 56
rect 5 6 9 56
<< polysilicon >>
rect 2 56 4 59
rect 2 -10 4 6
rect 2 -34 4 -30
<< polycontact >>
rect -2 -5 2 -1
<< metal1 >>
rect -9 61 16 64
rect -3 56 1 61
rect 5 -1 9 6
rect -9 -5 -2 -1
rect 5 -5 16 -1
rect 5 -10 9 -5
rect -3 -35 1 -30
rect -9 -38 16 -35
<< labels >>
rlabel metal1 3 -37 3 -37 1 gnd
rlabel metal1 -6 -3 -6 -3 3 input
rlabel metal1 11 -3 11 -3 7 output
rlabel metal1 -1 63 -1 63 5 vdd
<< end >>
