magic
tech scmos
timestamp 1613669700
<< nwell >>
rect 375 38 381 101
<< metal1 >>
rect 373 99 383 102
rect -19 33 0 37
rect 375 33 381 37
rect 401 33 418 37
rect -19 -33 -13 33
rect 375 2 381 3
rect 374 -3 406 2
rect 413 -33 418 33
rect -19 -37 1 -33
rect 372 -37 418 -33
use inverter  inverter_0
array 0 14 25 0 0 102
timestamp 1613668438
transform 1 0 9 0 1 38
box -9 -38 16 64
use inverter  inverter_2
timestamp 1613668438
transform 1 0 390 0 1 38
box -9 -38 16 64
use inverter  inverter_1
array 0 14 25 0 0 -102
timestamp 1613668438
transform 1 0 9 0 -1 -38
box -9 -38 16 64
<< labels >>
rlabel metal1 -2 35 -2 35 1 m1
rlabel space 25 35 25 35 1 m2
rlabel space 51 35 51 35 1 m3
rlabel space 76 35 76 35 1 m4
rlabel space 100 35 100 35 1 m5
rlabel space 125 35 125 35 1 m6
rlabel space 149 35 149 35 1 m7
rlabel space 176 36 176 36 1 m8
rlabel space 200 35 200 35 1 m9
rlabel space 224 35 224 35 1 m10
rlabel space 250 35 250 35 1 m11
rlabel space 275 34 275 34 1 m12
rlabel space 299 35 299 35 1 m13
rlabel space 325 36 325 36 1 m14
rlabel space 350 35 350 35 1 m15
rlabel metal1 376 35 376 35 1 m16
rlabel metal1 406 35 406 35 1 m17
rlabel space 350 -34 350 -34 1 m18
rlabel space 325 -35 325 -35 1 m19
rlabel space 297 -35 297 -35 1 m20
rlabel space 275 -35 275 -35 1 m21
rlabel space 248 -36 248 -36 1 m22
rlabel space 224 -35 224 -35 1 m23
rlabel space 199 -35 199 -35 1 m24
rlabel space 174 -35 174 -35 1 m25
rlabel space 150 -35 150 -35 1 m26
rlabel space 125 -35 125 -35 1 m27
rlabel space 100 -35 100 -35 1 m28
rlabel space 74 -35 74 -35 1 m29
rlabel space 49 -35 49 -35 1 m30
rlabel space 25 -36 25 -36 1 m31
<< end >>
