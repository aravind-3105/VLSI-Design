VLSI Assignment Question 7a
* Answers to question 7a
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.18u
.param W_N = 1.8u
.param width_P=20*LAMBDA
.param width_N=10*LAMBDA
.global gnd vdd

Vdd	 vdd gnd 'SUPPLY'
* Vin	 a	 gnd	0V
vin a 0 pulse 0 1.8 0ns 1ns 1ns 10ns 20ns

M1  b  a  vdd  vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2  b  a  gnd   gnd     CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M3  b  c  vdd   vdd     CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M4  b  c  gnd   gnd    CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

Cout c gnd 100f

.tran 0.1n 200n

.control
run
*plot v(a)
*plot v(b)
plot  v(c) v(a)

hardcopy fig_inv_trans.eps v(a) v(c)
.endc













