* SPICE3 file created from new.ext - technology: scmos

.option scale=0.09u

M1000 a_13_n25# a_6_n5# a_5_6# w_n1_0# pfet w=54 l=3
+  ad=270 pd=118 as=540 ps=236
M1001 a_38_n25# a_13_n25# a_5_6# w_n1_0# pfet w=54 l=3
+  ad=270 pd=118 as=0 ps=0
M1002 a_13_n25# a_6_n5# a_5_n25# Gnd nfet w=17 l=3
+  ad=85 pd=44 as=170 ps=88
M1003 a_38_n25# a_13_n25# a_5_n25# Gnd nfet w=17 l=3
+  ad=85 pd=44 as=0 ps=0
C0 w_n1_0# gnd! 3.4fF
