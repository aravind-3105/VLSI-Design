magic
tech scmos
timestamp 1613809452
<< metal1 >>
rect -18 68 360 72
rect -18 -68 -12 68
rect -9 28 7 32
rect 14 28 31 32
rect 38 28 54 32
rect 62 28 78 32
rect 86 28 102 32
rect 110 28 126 32
rect 134 28 150 32
rect 158 28 174 32
rect 182 28 198 32
rect 206 28 222 32
rect 230 28 246 32
rect 254 28 270 32
rect 278 28 294 32
rect 302 28 318 32
rect 326 28 342 32
rect 350 28 400 32
rect -9 -28 -3 28
rect 0 -4 384 4
rect 394 -28 400 28
rect -9 -32 6 -28
rect 17 -32 33 -28
rect 42 -32 58 -28
rect 66 -32 82 -28
rect 90 -32 106 -28
rect 114 -32 130 -28
rect 138 -32 154 -28
rect 162 -32 178 -28
rect 185 -32 201 -28
rect 210 -32 226 -28
rect 234 -32 250 -28
rect 258 -32 274 -28
rect 281 -32 297 -28
rect 305 -32 321 -28
rect 329 -32 345 -28
rect 353 -32 369 -28
rect 384 -32 400 -28
rect -18 -72 9 -68
use inverter_wo_label_Q5  inverter_wo_label_Q5_0
array 0 14 24 0 0 72
timestamp 1613681421
transform 1 0 0 0 1 33
box 0 -33 24 39
use inverter_wo_label_Q5  inverter_wo_label_Q5_1
array 0 15 -24 0 0 -72
timestamp 1613681421
transform -1 0 24 0 -1 -33
box 0 -33 24 39
<< labels >>
rlabel metal1 0 -4 384 4 1 gnd
rlabel metal1 0 68 360 72 5 vdd
rlabel metal1 -9 28 7 32 1 M1
rlabel metal1 14 28 31 32 1 M2
rlabel metal1 38 28 54 32 1 M3
rlabel metal1 62 28 78 32 1 M4
rlabel metal1 86 28 102 32 1 M5
rlabel metal1 110 28 126 32 1 M6
rlabel metal1 134 28 150 32 1 M7
rlabel metal1 158 28 174 32 1 M8
rlabel metal1 182 28 198 32 1 M9
rlabel metal1 206 28 222 32 1 M10
rlabel metal1 230 28 246 32 1 M11
rlabel metal1 254 28 270 32 1 M12
rlabel metal1 278 28 294 32 1 M13
rlabel metal1 302 28 318 32 1 M14
rlabel metal1 326 28 342 32 1 M15
rlabel metal1 350 28 366 32 1 M16
rlabel metal1 353 -32 369 -28 1 M17
rlabel metal1 329 -32 345 -28 1 M18
rlabel metal1 305 -32 321 -28 1 M19
rlabel metal1 281 -32 297 -28 1 M20
rlabel metal1 258 -32 274 -28 1 M21
rlabel metal1 234 -32 250 -28 1 M22
rlabel metal1 210 -32 226 -28 1 M23
rlabel metal1 185 -32 201 -28 1 M24
rlabel metal1 162 -32 178 -28 1 M25
rlabel metal1 138 -32 154 -28 1 M26
rlabel metal1 114 -32 130 -28 1 M27
rlabel metal1 90 -32 106 -28 1 M28
rlabel metal1 66 -32 82 -28 1 M29
rlabel metal1 42 -32 58 -28 1 M30
rlabel metal1 17 -32 33 -28 1 M31
<< end >>
