.param supply = 1.2V
.param length = 130n
.param wpmos=2500n wnmos=1000n

vsupply vdd 0 {supply}
vgnd vss 0 0V

Inputs to transistors
vin vgs vss dc 0

******************MOSFETs drain gate source body
Mpa vout vgs vdd vdd pmos l={length} w={wpmos} ; pmos
Mna vout vgs vss vss nmos l={length} w={wnmos} ; nmos

Cload vout vss1 200f
vdc0 vss1 vss dc 0V

.dc vin 0 1.2 0.1
*.tran 0.1n 500n 0 0.1n.
.save all @vsupply[p]

.control
run
plot v(vgs) v(vout)
.endc
.End