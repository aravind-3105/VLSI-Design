magic
tech scmos
timestamp 1613141391
<< nwell >>
rect 0 0 53 21
<< ntransistor >>
rect 11 -17 13 -13
rect 40 -17 42 -13
<< ptransistor >>
rect 11 7 13 15
rect 40 7 42 15
<< ndiffusion >>
rect 10 -17 11 -13
rect 13 -17 14 -13
rect 39 -17 40 -13
rect 42 -17 43 -13
<< pdiffusion >>
rect 10 7 11 15
rect 13 7 14 15
rect 39 7 40 15
rect 42 7 43 15
<< ndcontact >>
rect 6 -17 10 -13
rect 14 -17 18 -13
rect 35 -17 39 -13
rect 43 -17 47 -13
<< pdcontact >>
rect 6 7 10 15
rect 14 7 18 15
rect 35 7 39 15
rect 43 7 47 15
<< polysilicon >>
rect 11 15 13 18
rect 40 15 42 18
rect 11 -13 13 7
rect 40 -13 42 7
rect 11 -20 13 -17
rect 40 -20 42 -17
<< polycontact >>
rect 7 -7 11 -3
rect 36 -7 40 -3
<< metal1 >>
rect 0 20 53 25
rect 6 15 10 20
rect 35 15 39 20
rect 14 -3 18 7
rect 43 -3 47 7
rect -2 -7 7 -3
rect 14 -7 36 -3
rect 43 -7 56 -3
rect 14 -13 18 -7
rect 43 -13 47 -7
rect 6 -23 10 -17
rect 35 -23 39 -17
rect 6 -27 47 -23
<< labels >>
rlabel metal1 -1 -5 -1 -5 3 in
rlabel metal1 27 -5 27 -5 1 mid
rlabel metal1 54 -5 54 -5 7 out
rlabel metal1 24 23 24 23 5 vdd
rlabel metal1 26 -25 26 -25 1 gnd
<< end >>
