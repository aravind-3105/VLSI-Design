magic
tech scmos
timestamp 1613133646
<< nwell >>
rect 0 0 25 23
<< ntransistor >>
rect 11 -13 13 -9
<< ptransistor >>
rect 11 6 13 14
<< ndiffusion >>
rect 10 -13 11 -9
rect 13 -13 14 -9
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
<< ndcontact >>
rect 6 -13 10 -9
rect 14 -13 18 -9
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
<< polysilicon >>
rect 11 14 13 17
rect 11 -9 13 6
rect 11 -18 13 -13
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 0 19 25 28
rect 6 14 10 19
rect 14 -1 18 6
rect -6 -5 7 -1
rect 14 -5 31 -1
rect 14 -9 18 -5
rect 6 -20 10 -13
rect -2 -26 22 -20
<< labels >>
rlabel metal1 7 -24 7 -24 1 gnd
rlabel pdcontact 8 10 8 10 1 Psrc
rlabel pdcontact 16 10 16 10 1 Pdrn
rlabel metal1 -3 -3 -3 -3 3 input
rlabel metal1 27 -3 27 -3 7 output
rlabel ndcontact 8 -11 8 -11 1 Nsrc
rlabel ndcontact 16 -11 16 -11 1 Ndrn
rlabel metal1 9 24 9 24 5 Vdd
<< end >>
