magic
tech scmos
timestamp 1617455408
<< nwell >>
rect 0 0 24 26
<< ntransistor >>
rect 11 -14 13 -8
<< ptransistor >>
rect 11 6 13 18
<< ndiffusion >>
rect 10 -14 11 -8
rect 13 -14 14 -8
<< pdiffusion >>
rect 10 6 11 18
rect 13 6 14 18
<< ndcontact >>
rect 6 -14 10 -8
rect 14 -14 18 -8
<< pdcontact >>
rect 6 6 10 18
rect 14 6 18 18
<< polysilicon >>
rect 11 18 13 21
rect 11 -8 13 6
rect 11 -17 13 -14
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 0 23 24 26
rect 6 18 10 23
rect 14 -1 18 6
rect 0 -5 7 -1
rect 14 -5 24 -1
rect 14 -8 18 -5
rect 6 -18 10 -14
rect 0 -21 24 -18
<< labels >>
rlabel metal1 4 -3 4 -3 3 inp
rlabel metal1 18 -3 18 -3 1 out
rlabel metal1 7 -19 7 -19 1 gnd
rlabel metal1 8 24 8 24 5 vdd
<< end >>
