* SPICE3 file created from double_inverter.ext - technology: scmos
* Answers to question 3
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.option scale=0.09u
.global gnd vdd

Vdd vdd gnd 1.8V
vin in 0 0V 

M1000 mid in vdd w_0_0# CMOSP w=50 l=2
+  ad=250 pd=110 as=500 ps=220

M1001 out mid vdd w_0_0# CMOSP w=50 l=2
+  ad=250 pd=110 as=0 ps=0

M1002 mid in gnd gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100

M1003 out mid gnd gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0

C0 w_0_0# gnd 2.9fF

.dc vin 0 1.8 0.01

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
let a = v(mid)
let b = deriv(v(mid))/deriv(v(in))
let c= 1V
set curplottitle="AravindNarayanan-2019102014-Q3d-VTC"
plot  a c
set curplottitle="AravindNarayanan-2019102014-Q3d-SLOPE"
plot  b c

hardcopy fig_Q3d.eps v(mid) deriv(v(mid))/deriv(v(in)) c
.endc


