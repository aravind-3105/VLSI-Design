
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.global gnd vdd

Vdd	vg	gnd	'SUPPLY'
VGS G gnd 1.8V



M1 G vin vc gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

Cout vc gnd 100f

.dc VGS 0 1.8 0.01


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
let x = (-vout#branch)
set curplottitle="Id vs Vgs Characteristics"
plot x 

hardcopy fig_inv_trans.eps (-vout#branch)
.endc
