VLSI Assignment Question 3ii
* Answers to question 3ii
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_P={20*LAMBDA}
.global gnd vdd

VGS G gnd 0
VDS D gnd 1.8V
VBS B D 900mV

M1 D G gnd B CMOSP W={width_P} L={2*LAMBDA} 
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+ AD={5*width_P*LAMBDA}

.dc VGS 0 1.8 0.001


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
let x = (-VDS#branch)
set curplottitle="Id vs Vgs Characteristics"
plot x 

let y = sqrt(-VDS#branch)
set curplottitle="sqrt(Id) vs Vgs Characteristics"
plot y

let z = deriv(sqrt(-VDS#branch))/deriv(V(G))
set curplottitle="First derivative Characteristics"
plot z

hardcopy fig_Q3iiPMOS.eps (-VDS#branch) sqrt(-VDS#branch) deriv(sqrt(-VDS#branch))/deriv(V(G))
.endc
