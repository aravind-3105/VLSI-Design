VLSI Assignment Question 3i
* Answers to question 3i
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.global gnd vdd

VGS G gnd 0V
VDS D gnd 1.8V
VBS B gnd 0V

M1 D G gnd B CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA}

.dc VGS 0 1.8 0.01


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
let x = (-VDS#branch)
let y = sqrt(-VDS#branch)
let z = deriv(sqrt(-VDS#branch))
let zz = deriv(sqrt(-VDS#branch))/deriv(V(G))

set curplottitle="Id vs Vgs Characteristics"
plot x 

set curplottitle="deriv(Id) vs Vgs Characteristics"
plot y

set curplottitle="Id vs Vgs Characteristics"
plot z

hardcopy fig_Q3iNMOS.eps (-VDS#branch)
.endc
