* SPICE3 file created from ring.ext - technology: scmos

.option scale=0.09u

M1000 inverter_1[0]/a_4_n30# m1 inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=3750 ps=1650
M1001 inverter_1[0]/a_4_n30# m1 inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=3100 ps=1550
M1002 inverter_1[1]/a_4_n30# inverter_1[0]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1003 inverter_1[1]/a_4_n30# inverter_1[0]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 inverter_1[2]/a_4_n30# inverter_1[1]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1005 inverter_1[2]/a_4_n30# inverter_1[1]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 inverter_1[3]/a_4_n30# inverter_1[2]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1007 inverter_1[3]/a_4_n30# inverter_1[2]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1008 inverter_1[4]/a_4_n30# inverter_1[3]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1009 inverter_1[4]/a_4_n30# inverter_1[3]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 inverter_1[5]/a_4_n30# inverter_1[4]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1011 inverter_1[5]/a_4_n30# inverter_1[4]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1012 inverter_1[6]/a_4_n30# inverter_1[5]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1013 inverter_1[6]/a_4_n30# inverter_1[5]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1014 inverter_1[7]/a_4_n30# inverter_1[6]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1015 inverter_1[7]/a_4_n30# inverter_1[6]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1016 inverter_1[8]/a_4_n30# inverter_1[7]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1017 inverter_1[8]/a_4_n30# inverter_1[7]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1018 inverter_1[9]/a_4_n30# inverter_1[8]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1019 inverter_1[9]/a_4_n30# inverter_1[8]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1020 inverter_1[10]/a_4_n30# inverter_1[9]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1021 inverter_1[10]/a_4_n30# inverter_1[9]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1022 inverter_1[11]/a_4_n30# inverter_1[10]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1023 inverter_1[11]/a_4_n30# inverter_1[10]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1024 inverter_1[12]/a_4_n30# inverter_1[11]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1025 inverter_1[12]/a_4_n30# inverter_1[11]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1026 inverter_1[13]/a_4_n30# inverter_1[12]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1027 inverter_1[13]/a_4_n30# inverter_1[12]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1028 m17 inverter_1[13]/a_4_n30# inverter_1[0]/vdd inverter_1[0]/w_n9_0# pfet w=50 l=2
+  ad=500 pd=220 as=0 ps=0
M1029 m17 inverter_1[13]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1030 m17 m16 inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=0 pd=0 as=4000 ps=1760
M1031 m17 m16 inverter_2/gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 inverter_0[0]/a_4_n30# m1 inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1033 inverter_0[0]/a_4_n30# m1 inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1034 inverter_0[1]/a_4_n30# inverter_0[0]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1035 inverter_0[1]/a_4_n30# inverter_0[0]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1036 inverter_0[2]/a_4_n30# inverter_0[1]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1037 inverter_0[2]/a_4_n30# inverter_0[1]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1038 inverter_0[3]/a_4_n30# inverter_0[2]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1039 inverter_0[3]/a_4_n30# inverter_0[2]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1040 inverter_0[4]/a_4_n30# inverter_0[3]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1041 inverter_0[4]/a_4_n30# inverter_0[3]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1042 inverter_0[5]/a_4_n30# inverter_0[4]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1043 inverter_0[5]/a_4_n30# inverter_0[4]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1044 inverter_0[6]/a_4_n30# inverter_0[5]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1045 inverter_0[6]/a_4_n30# inverter_0[5]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1046 inverter_0[7]/a_4_n30# inverter_0[6]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1047 inverter_0[7]/a_4_n30# inverter_0[6]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1048 inverter_0[8]/a_4_n30# inverter_0[7]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1049 inverter_0[8]/a_4_n30# inverter_0[7]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1050 inverter_0[9]/a_4_n30# inverter_0[8]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1051 inverter_0[9]/a_4_n30# inverter_0[8]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1052 inverter_0[10]/a_4_n30# inverter_0[9]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1053 inverter_0[10]/a_4_n30# inverter_0[9]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1054 inverter_0[11]/a_4_n30# inverter_0[10]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1055 inverter_0[11]/a_4_n30# inverter_0[10]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1056 inverter_0[12]/a_4_n30# inverter_0[11]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1057 inverter_0[12]/a_4_n30# inverter_0[11]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1058 inverter_0[13]/a_4_n30# inverter_0[12]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1059 inverter_0[13]/a_4_n30# inverter_0[12]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1060 m16 inverter_0[13]/a_4_n30# inverter_2/vdd w_375_38# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1061 m16 inverter_0[13]/a_4_n30# inverter_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 inverter_1[0]/vdd inverter_1[0]/w_n9_0# 1.6fF
C1 inverter_2/vdd w_375_38# 1.7fF
C2 inverter_2/gnd gnd! 3.0fF
C3 w_375_38# gnd! 26.1fF
C4 inverter_1[0]/w_n9_0# gnd! 23.7fF
