VLSI Assignment Question 3S=a
* Answers to question 3a
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N=20*LAMBDA
.param width_P=2.5*width_N
.global gnd vdd

Vdd vdd gnd 1.8V
vin x 0 0V 

M1      y       x       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2      y       x       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M3      z       y       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M4      z       y       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

Cout z gnd 100f

.dc vin 0 1.8 0.0001



.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
let a = v(y)
let b = deriv(v(y))/deriv(v(x))
set curplottitle="AravindNarayanan-2019102014-Q3a-VTC"
plot  a
set curplottitle="AravindNarayanan-2019102014-Q3a-SLOPE"
plot  b

hardcopy fig_Q3a.eps v(z) deriv(v(y))/deriv(v(x))
.endc





