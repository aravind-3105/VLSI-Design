.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 'SUPPLY'
vin input gnd pulse 0 1.8 0ns 1ns 1ns 10ns 20ns


M1000 output input Vdd w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=125 ps=60
M1001 output input gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 w_0_0# gnd 1.1fF

.tran 0.01n 200n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
set curplottitle="v(out)"
plot v(input) v(output)
hardcopy WithLabel.eps v(input) v(output)
.endc

.end