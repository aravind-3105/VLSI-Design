* SPICE3 file created from oscillator.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

M1000 m2 m1 vdd vdd CMOSP w=50 l=2
+  ad=250 pd=110 as=750 ps=330
M1001 m2 m1 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=300 ps=150

M1002 m3 m2 vdd vdd CMOSP w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1003 m3 m2 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0

M1004 m1 m3 vdd vdd CMOSP w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1005 m1 m3 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 vdd gnd 4.7fF

.ic v(m1) = 'SUPPLY'
.tran 0.001n 2n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
set curplottitle="v(out)"
plot v(m1) v(m2) v(m3)
hardcopy RIng_3.eps v(m1) v(m2) v(m3)
.endc