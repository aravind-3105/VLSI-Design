magic
tech scmos
timestamp 1613517333
<< nwell >>
rect -1 0 49 68
<< ntransistor >>
rect 10 -25 13 -8
rect 35 -25 38 -8
<< ptransistor >>
rect 10 6 13 60
rect 35 6 38 60
<< ndiffusion >>
rect 9 -25 10 -8
rect 13 -25 14 -8
rect 34 -25 35 -8
rect 38 -25 39 -8
<< pdiffusion >>
rect 9 6 10 60
rect 13 6 14 60
rect 34 6 35 60
rect 38 6 39 60
<< ndcontact >>
rect 5 -25 9 -8
rect 14 -25 18 -8
rect 30 -25 34 -8
rect 39 -25 43 -8
<< pdcontact >>
rect 5 6 9 60
rect 14 6 18 60
rect 30 6 34 60
rect 39 6 43 60
<< polysilicon >>
rect 10 60 13 63
rect 35 60 38 63
rect 10 -8 13 6
rect 35 -8 38 6
rect 10 -32 13 -25
rect 35 -32 38 -25
<< polycontact >>
rect 6 -5 10 -1
rect 31 -5 35 -1
<< metal1 >>
rect -1 65 49 68
rect 5 60 9 65
rect 30 60 34 65
rect 14 -1 18 6
rect 39 -1 43 6
rect -6 -5 6 -1
rect 14 -5 31 -1
rect 39 -5 57 -1
rect 14 -8 18 -5
rect 39 -8 43 -5
rect 5 -34 9 -25
rect 30 -34 34 -25
rect 5 -37 43 -34
<< labels >>
rlabel metal1 1 -3 1 -3 1 in
rlabel metal1 25 -3 25 -3 1 x
rlabel metal1 51 -3 51 -3 1 out
rlabel metal1 25 67 25 67 5 vdd
rlabel metal1 17 -36 17 -36 1 gnd
<< end >>
