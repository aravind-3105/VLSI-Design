* SPICE3 file created from optimized_ring_oscillator.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 'SUPPLY'

M1000 M2 M1 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1001 M2 M1 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1002 M3 M2 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1003 M3 M2 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1004 M4 M3 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1005 M4 M3 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1006 M5 M4 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1007 M5 M4 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1008 M6 M5 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1009 M6 M5 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1010 M7 M6 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1011 M7 M6 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1012 M8 M7 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1013 M8 M7 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1014 M9 M8 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1015 M9 M8 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1016 M10 M9 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1017 M10 M9 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1018 M11 M10 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1019 M11 M10 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1020 M12 M11 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1021 M12 M11 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1022 M13 M12 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1023 M13 M12 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1024 M14 M13 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1025 M14 M13 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1026 M15 M14 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1027 M15 M14 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1028 M16 M15 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1029 M16 M15 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1030 M17 M16 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1031 M17 M16 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1032 M18 M17 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1033 M18 M17 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1034 M19 M18 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1035 M19 M18 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1036 M20 M19 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1037 M20 M19 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1038 M21 M20 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1039 M21 M20 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1040 M22 M21 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1041 M22 M21 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1042 M23 M22 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1043 M23 M22 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1044 M24 M23 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1045 M24 M23 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1046 M25 M24 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1047 M25 M24 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1048 M26 M25 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1049 M26 M25 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1050 M27 M26 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1051 M27 M26 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1052 M28 M27 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1053 M28 M27 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1054 M29 M28 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1055 M29 M28 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1056 M30 M29 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1057 M30 M29 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1058 M31 M30 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1059 M31 M30 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

M1060 M1 M31 vdd vdd CMOSP w=25 l=2
+  ad=125 pd=60 as=3875 ps=1860
M1061 M1 M31 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=1550 ps=930



C0 vdd vdd 1.2fF
C1 vdd vdd 1.2fF
C2 vdd gnd 2.3fF
C3 vdd gnd 13.4fF
C4 gnd gnd 3.2fF
C5 M16 gnd 1.0fF
C6 vdd gnd 14.3fF
C7 M30 gnd 1.1fF
C8 M31 gnd 1.2fF
C9 M1 gnd 2.1fF

.ic v(M1) = 'SUPPLY'
.tran 1n 20n

** MEASURING DELAYS
.measure tran tpdr
+ TRIG v(M1) VAL='SUPPLY/2' FALL=1
+ TARG v(M2) VAL='SUPPLY/2' RISE=1

.measure tran tpdf
+ TRIG v(M1) VAL='SUPPLY/2' RISE=1
+ TARG v(M2) VAL='SUPPLY/2' FALL=1

.measure tran tpd param='(tpdr+tpdf)/2' goal=0


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
set curplottitle="AravindNarayanan-2019102014-Q5-b(i)-Optimized"
plot v(M1)
hardcopy Optimized_Ring_Oscillator.eps v(M1)
.endc

.end
