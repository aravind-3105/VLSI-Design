.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={2.5*width_N}
.global gnd vdd

.option scale=0.09u

M1000 17 16 vdd basicinv_0[0]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=3875 ps=1860
M1001 17 16 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=1550 ps=930
M1002 18 17 vdd basicinv_0[1]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1003 18 17 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1004 19 18 vdd basicinv_0[2]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1005 19 18 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1006 20 19 vdd basicinv_0[3]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1007 20 19 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1008 21 20 vdd basicinv_0[4]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1009 21 20 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1010 22 21 vdd basicinv_0[5]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1011 22 21 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1012 23 22 vdd basicinv_0[6]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1013 23 22 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1014 24 23 vdd basicinv_0[7]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1015 24 23 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1016 25 24 vdd basicinv_0[8]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1017 25 24 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1018 26 25 vdd basicinv_0[9]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1019 26 25 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1020 27 26 vdd basicinv_0[10]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1021 27 26 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1022 28 27 vdd basicinv_0[11]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1023 28 27 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1024 29 28 vdd basicinv_0[12]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1025 29 28 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 30 29 vdd basicinv_0[13]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1027 30 29 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1028 in 30 vdd basicinv_0[14]/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1029 in 30 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1030 16 15 vdd basicinv_1/w_0_0# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1031 16 15 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1032 15 14 vdd w_2_423# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1033 15 14 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1034 14 13 vdd w_2_393# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1035 14 13 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1036 13 12 vdd w_2_363# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1037 13 12 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1038 12 11 vdd w_2_333# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1039 12 11 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 11 10 vdd w_2_303# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1041 11 10 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1042 10 9 vdd w_2_273# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1043 10 9 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1044 9 8 vdd w_2_243# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1045 9 8 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1046 8 7 vdd w_2_213# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1047 8 7 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1048 7 6 vdd w_2_183# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1049 7 6 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 6 5 vdd w_2_153# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1051 6 5 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1052 5 4 vdd w_2_123# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1053 5 4 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1054 4 3 vdd w_2_93# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1055 4 3 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1056 3 2 vdd w_2_63# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1057 3 2 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1058 2 1 vdd w_2_33# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1059 2 1 gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 1 in vdd w_2_3# CMOSP w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1061 1 in gnd gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0

C0 w_2_33# gnd 1.0fF
C1 w_2_63# gnd 1.0fF
C2 w_2_93# gnd 1.0fF
C3 w_2_123# gnd 1.0fF
C4 w_2_153# gnd 1.0fF
C5 w_2_183# gnd 1.0fF
C6 w_2_213# gnd 1.0fF
C7 w_2_243# gnd 1.0fF
C8 w_2_273# gnd 1.0fF
C9 w_2_303# gnd 1.0fF
C10 w_2_333# gnd 1.0fF
C11 w_2_363# gnd 1.0fF
C12 w_2_393# gnd 1.0fF
C13 w_2_423# gnd 1.0fF
C14 gnd gnd 6.4fF
C15 basicinv_1/w_0_0# gnd 1.0fF
C16 vdd gnd 8.4fF

Vdd	vdd	gnd	'SUPPLY'

.ic v(in) = 'SUPPLY'
.tran 1n 100n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))

run
set curplottitle="v(in)"
plot v(in)

.endc