VLSI Assignment Question 5
* Answers to question 5
.include TSMC_180nm.txt
.param SUPPLY=1.8V
.param LAMBDA=0.09u
.param width_N=10*LAMBDA
.param width_P=2.5*width_N
.global gnd vdd

Vdd vdd gnd 1.8V
vin in gnd pulse 0 1.8 0ns 0ns 0ns 10ns 20ns


M1      out       in       gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2      out       in       vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}


*.ic v(in)= 1.8V
.tran 0.01n 50n



** MEASURING DELAYS
.measure tran tpdr
+ TRIG v(in) VAL='SUPPLY/2' FALL=1
+ TARG v(out) VAL='SUPPLY/2' RISE=1

.measure tran tpdf
+ TRIG v(in) VAL='SUPPLY/2' RISE=1
+ TARG v(out) VAL='SUPPLY/2' FALL=1

.measure tran tpd param='(tpdr+tpdf)/2' goal=0


.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
*plot v(a)
*plot v(b)
set curplottitle="AravindNarayanan-2019102014-Q5-a"
plot  v(in) v(out)

hardcopy fig_Q5a_single.eps v(in) v(out)
.endc

